library verilog;
use verilog.vl_types.all;
entity BK_adder_t is
end BK_adder_t;
